module porta_not_behav(a, y);
  input a;
  output y;
  assign y = ~a;
endmodule