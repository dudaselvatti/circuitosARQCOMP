module porta_xor_behav(a, b, y);
    input a, b;
    output y;
    assign y = a ^ b;
endmodule