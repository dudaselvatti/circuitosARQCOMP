module porta_or_behav(a, b, y);
  input a, b;
  output y;
  assign y = a | b;
endmodule